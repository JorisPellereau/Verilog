module wait_duration #(
		       )
   ();

   wait_duration_intf wait_duration_if();
   
endmodule // wait_duration
