interface master_axi4lite_intf #(parameter G_AXI4LITE_ADDR_WIDTH = 32,
				 parameter G_AXI4LITE_DATA_WIDTH = 32
				 );

endinterface // master_axi4lite_intf
