//                              -*- Mode: Verilog -*-
// Filename        : testbench_class.sv
// Description     : Testbench class
// Author          : JorisP
// Created On      : Sat May  1 20:40:14 2021
// Last Modified By: JorisP
// Last Modified On: Sat May  1 20:40:14 2021
// Update Count    : 0
// Status          : Unknown, Use with caution!

`include "tb_tasks.sv"

class testbench_class;

   // == STATIC Functions ==

   
   
   // ======================
endclass // testbench_class
