interface wait_duration_intf; 
   
   logic clk;
        
endinterface // wait_duration_intf

