//                              -*- Mode: Verilog -*-
// Filename        : tb_interfaces.sv
// Description     : TB Interfaces
// Author          : JorisP
// Created On      : Fri Nov 13 19:49:50 2020
// Last Modified By: JorisP
// Last Modified On: Fri Nov 13 19:49:50 2020
// Update Count    : 0
// Status          : Unknown, Use with caution!

// == INTERFACES ==
  /* interface wait_event_intf #(
     parameter WAIT_SIZE  = 5,
     parameter WAIT_WIDTH = 1
   );
   
   logic wait_en;   
   logic sel_wtr_wtf;
   logic [31:0] max_timeout;
   logic [WAIT_WIDTH - 1 : 0] wait_signals [WAIT_SIZE];   
   logic 	wait_done;
   
   endinterface*/ // wait_event_int
   
   // ===============
