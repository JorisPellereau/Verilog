module tb_test

endmodule // tb_test
