/*
 *
 *  interface.sv
 * 
 */

interface intf (input logic clk, rst_n);
   logic i_en_cnt;   
   
endinterface //

