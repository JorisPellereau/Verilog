jorisp@jorisp-VirtualBox.2920:1619630158